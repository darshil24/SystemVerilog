
//Greg Stitt
//University of Florida
‘timescale 1ns / 10ps
/* the software tool is instructed to use time units of 1 nanosecond,
and a precision of 10 picoseconds, which is 2 decimal places, relative to 1 nanosecond. */