//Greg Stitt
//University of Florida


module add(in1, in2,sum,carry);	
		parameter WIDTH = 8;
		input    in1 [WIDTH-1 : 0];
		input    in2 [WIDTH-1 : 0];
		input  	 sum[WIDTH-1 : 0];
		output   carry;
		logic  	 carry;
		logic 	 sum;
	
always  @(in1, in2)
	
endmodule



















